// Copyright 2023 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Authors:
// - Thomas Benz <tbenz@iis.ee.ethz.ch>
// - Paul Scheffler <paulsc@iis.ee.ethz.ch>
//
// Based on work of:
// - Fabian Schuiki <fschuiki@iis.ee.ethz.ch>
// - Florian Zaruba <zarubaf@iis.ee.ethz.ch>
//
// Automatically generated by gen_model.py

module delay_line_D4_O1_6P000 (
    input  logic       clk_i,
    input  logic [3:0] delay_i,
    output logic [0:0] clk_o
);

    assign #(real'(delay_i) * 0.4ns/6.000 + 0.3ns) clk_o[0] = clk_i;

endmodule

